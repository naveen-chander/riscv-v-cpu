add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM1/inst/wea[0]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM2/inst/wea[0]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM3/inst/wea[0]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM4/inst/wea[0]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM5/inst/wea[0]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM6/inst/wea[0]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/DMEM7/inst/wea[0]}} 


add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(0)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(1)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(2)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(3)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(4)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(5)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(6)\/vrf_gen/vec_reg[28]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(7)\/vrf_gen/vec_reg[28]}}


add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(1)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(0)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(2)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(3)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(4)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(5)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(6)\/vrf_gen/vec_reg[29]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(7)\/vrf_gen/vec_reg[29]}}

add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(0)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(1)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(2)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(3)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(4)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(5)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(6)\/vrf_gen/vec_reg[30]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(7)\/vrf_gen/vec_reg[30]}}

add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(0)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(1)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(2)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(3)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(4)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(5)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(6)\/vrf_gen/vec_reg[31]}} 
add_wave {{/FPGA_WRAPPER_TEST/FW1/cpu1/fdem/Pipeline/VECTOR_UNIT/VEC_EXE_UNIT/wrapper_vhd/VECTOR_EXE_UNIT_PIPE/\GEN_VRFS(7)\/vrf_gen/vec_reg[31]}}


